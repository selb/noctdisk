# edlin.sv - messages file (Swedish version)
# 
# Author: Gregory Pietsch
# 
# DESCRIPTION:
# 
# This file contains #defines for all the message strings in edlin.
# For internationalization fun, just translate the messages in this
# file.
# 
# The strings were generated using ESR's cstrings program and moved
# here.
# 
# 
# 
1.0:Jj
1.1: :  \b
1.2:O.K.?  \b
1.3:Intrade misstag.
1.4:%s: %lu lina l�ste\n
1.5:%s: %lu linjen l�ste\n
1.6:%s: %lu lina var skrev\n
1.7:%s: %lu linjen var skrev\n
1.8:%lu:%c%s\n
1.9:Pressa g� in till forts�tta
1.10:%lu:  \b
1.11:Inte grunda
1.12:%lu: %s\n
1.13:\nedlin has the following subcommands:\n
1.14:#                 redigera en enkel lina  [#],[#],#m        flytta
1.15:a                 till�gga                [#][,#]p          engelsk mynt sida
1.16:[#],[#],#,[#]c    kopia                   q                 l�mna
1.17:[#][,#]d          stryka                  [#][,#][?]r$,$    s�tta tillbaka
1.18:e<>               skriva & l�mna          [#][,#][?]s$      s�ka
1.19:[#]i              s�tta in                [#]t<>            l�ste
1.20:[#][,#]l          lista                   [#]w<>            skriva\n
1.21:var $ �ver �r en sn�re , <> �r en arkivnamnen,
1.22:# �r et antal (vilken Maj bli.current= lina, $=sist lina,
1.23:eller endera antal + eller - en annan antal).\n
1.24:, copyright (c) 2003 Gregory Pietsch
1.25:Den h�r program kommer med ABSOLUT INGEN GARANTIEN.
1.26:Den er fri mjukvaran, och du er v�lkommen till oml�gga den
1.27:under termen om GNU General Allm�nhet Licens endera version 2
1.28:om licens, eller, p� din valen, n�gon senare
1.29:version.\n
1.30:Ute om minne
1.31:Sn�re l�ngd misstag
1.32:Sn�re position misstag
1.33:Sjukling f�rbrukaren insatsen, anv�nda ? f�r hj�lp.
1.34:Nej arkivnamnen
1.35:Buffert alltf�r stor
1.36:Sjukling buffert position
1.37:MISSTAG: %s\n

# END OF FILE
